library verilog;
use verilog.vl_types.all;
entity test5_vlg_vec_tst is
end test5_vlg_vec_tst;
