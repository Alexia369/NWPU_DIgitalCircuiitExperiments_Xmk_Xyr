LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY XOR4_1 IS
PORT(A,B:IN STD_LOGIC;C:OUT STD_LOGIC);
END XOR4_1;
ARCHITECTURE fwm OF XOR4_1 IS
BEGIN
C<=A XOR B;
END;