library verilog;
use verilog.vl_types.all;
entity COUNT4_3_vlg_vec_tst is
end COUNT4_3_vlg_vec_tst;
