library verilog;
use verilog.vl_types.all;
entity iddisplay_1_vlg_vec_tst is
end iddisplay_1_vlg_vec_tst;
