library verilog;
use verilog.vl_types.all;
entity XOR4_1 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : out    vl_logic
    );
end XOR4_1;
