library verilog;
use verilog.vl_types.all;
entity iddisplay_1_vlg_check_tst is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        E               : in     vl_logic;
        F               : in     vl_logic;
        G               : in     vl_logic;
        H1              : in     vl_logic;
        H2              : in     vl_logic;
        H3              : in     vl_logic;
        H4              : in     vl_logic;
        L1              : in     vl_logic;
        L2              : in     vl_logic;
        L3              : in     vl_logic;
        L4              : in     vl_logic;
        OutCLK          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end iddisplay_1_vlg_check_tst;
