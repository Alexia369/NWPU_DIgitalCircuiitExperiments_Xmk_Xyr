library verilog;
use verilog.vl_types.all;
entity \32\ is
    port(
        D               : out    vl_logic_vector(6 downto 0);
        clk             : in     vl_logic
    );
end \32\;
