library verilog;
use verilog.vl_types.all;
entity DIVIDE4_4_vlg_check_tst is
    port(
        clk_out1        : in     vl_logic;
        clk_out2        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end DIVIDE4_4_vlg_check_tst;
