library verilog;
use verilog.vl_types.all;
entity iddisplay_1 is
    port(
        A               : out    vl_logic;
        clk             : in     vl_logic;
        B               : out    vl_logic;
        C               : out    vl_logic;
        D               : out    vl_logic;
        E               : out    vl_logic;
        F               : out    vl_logic;
        G               : out    vl_logic;
        H1              : out    vl_logic;
        H2              : out    vl_logic;
        H3              : out    vl_logic;
        H4              : out    vl_logic;
        L4              : out    vl_logic;
        L3              : out    vl_logic;
        L2              : out    vl_logic;
        L1              : out    vl_logic
    );
end iddisplay_1;
