library verilog;
use verilog.vl_types.all;
entity XOR4_1_vlg_vec_tst is
end XOR4_1_vlg_vec_tst;
