library verilog;
use verilog.vl_types.all;
entity test4_vlg_vec_tst is
end test4_vlg_vec_tst;
