library verilog;
use verilog.vl_types.all;
entity DIVIDE4_4_vlg_vec_tst is
end DIVIDE4_4_vlg_vec_tst;
