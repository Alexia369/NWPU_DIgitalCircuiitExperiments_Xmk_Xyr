library verilog;
use verilog.vl_types.all;
entity sdsy_vlg_vec_tst is
end sdsy_vlg_vec_tst;
