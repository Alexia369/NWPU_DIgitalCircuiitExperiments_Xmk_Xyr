library verilog;
use verilog.vl_types.all;
entity FINAL4_5_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        Switch          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end FINAL4_5_vlg_sample_tst;
