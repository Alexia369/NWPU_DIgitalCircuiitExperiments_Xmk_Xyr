library verilog;
use verilog.vl_types.all;
entity ROMuse_vlg_vec_tst is
end ROMuse_vlg_vec_tst;
