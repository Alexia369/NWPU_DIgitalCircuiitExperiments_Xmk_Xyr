library verilog;
use verilog.vl_types.all;
entity FINAL4_5_vlg_vec_tst is
end FINAL4_5_vlg_vec_tst;
