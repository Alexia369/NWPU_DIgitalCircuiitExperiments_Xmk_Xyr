library verilog;
use verilog.vl_types.all;
entity XOR4_1_vlg_check_tst is
    port(
        C               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end XOR4_1_vlg_check_tst;
