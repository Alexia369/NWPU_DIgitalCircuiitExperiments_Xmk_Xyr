library verilog;
use verilog.vl_types.all;
entity iddisplay_1_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end iddisplay_1_vlg_sample_tst;
