library verilog;
use verilog.vl_types.all;
entity FINAL4_5_vlg_check_tst is
    port(
        led             : in     vl_logic_vector(6 downto 0);
        sampler_rx      : in     vl_logic
    );
end FINAL4_5_vlg_check_tst;
